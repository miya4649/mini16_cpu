module default_code_mem
  #(
    parameter DATA_WIDTH=16,
    parameter ADDR_WIDTH=8
    )
  (
   input                         clk,
   input [(ADDR_WIDTH-1):0]      addr_r,
   input [(ADDR_WIDTH-1):0]      addr_w,
   input [(DATA_WIDTH-1):0]      data_in,
   input                         we,
   output reg [(DATA_WIDTH-1):0] data_out
   );

  reg [DATA_WIDTH-1:0]           ram [0:(1 << ADDR_WIDTH)-1];

  always @(posedge clk)
    begin
      data_out <= ram[addr_r];
      if (we)
        begin
          ram[addr_w] <= data_in;
        end
    end

  initial
    begin
      ram[16'h0000] = 16'h0000;
      ram[16'h0001] = 16'h2011;
      ram[16'h0002] = 16'h0000;
      ram[16'h0003] = 16'h0000;
      ram[16'h0004] = 16'h0000;
      ram[16'h0005] = 16'h0000;
      ram[16'h0006] = 16'h0000;
      ram[16'h0007] = 16'h2050;
      ram[16'h0008] = 16'h03b1;
      ram[16'h0009] = 16'h0000;
      ram[16'h000a] = 16'h0000;
      ram[16'h000b] = 16'h0000;
      ram[16'h000c] = 16'h0000;
      ram[16'h000d] = 16'h0000;
      ram[16'h000e] = 16'h2850;
      ram[16'h000f] = 16'h0471;
      ram[16'h0010] = 16'h0000;
      ram[16'h0011] = 16'h0000;
      ram[16'h0012] = 16'h0000;
      ram[16'h0013] = 16'h0000;
      ram[16'h0014] = 16'h0000;
      ram[16'h0015] = 16'h3050;
      ram[16'h0016] = 16'h2011;
      ram[16'h0017] = 16'h1ff0;
      ram[16'h0018] = 16'h3830;
      ram[16'h0019] = 16'h0000;
      ram[16'h001a] = 16'h0000;
      ram[16'h001b] = 16'h0000;
      ram[16'h001c] = 16'h2050;
      ram[16'h001d] = 16'h10d0;
      ram[16'h001e] = 16'h0000;
      ram[16'h001f] = 16'h0000;
      ram[16'h0020] = 16'h0000;
      ram[16'h0021] = 16'h0000;
      ram[16'h0022] = 16'h0000;
      ram[16'h0023] = 16'h009c;
      ram[16'h0024] = 16'h1069;
      ram[16'h0025] = 16'h0000;
      ram[16'h0026] = 16'h0000;
      ram[16'h0027] = 16'h0000;
      ram[16'h0028] = 16'h0000;
      ram[16'h0029] = 16'h0185;
      ram[16'h002a] = 16'h0000;
      ram[16'h002b] = 16'h0000;
      ram[16'h002c] = 16'h0000;
      ram[16'h002d] = 16'h0000;
      ram[16'h002e] = 16'h0000;
      ram[16'h002f] = 16'h21c1;
      ram[16'h0030] = 16'h3868;
      ram[16'h0031] = 16'h0144;
      ram[16'h0032] = 16'h0000;
      ram[16'h0033] = 16'h0000;
      ram[16'h0034] = 16'h0000;
      ram[16'h0035] = 16'h0000;
      ram[16'h0036] = 16'h0000;
      ram[16'h0037] = 16'h0000;
      ram[16'h0038] = 16'h0000;
      ram[16'h0039] = 16'h0000;
      ram[16'h003a] = 16'h0000;
      ram[16'h003b] = 16'h0000;
      ram[16'h003c] = 16'h0000;
      ram[16'h003d] = 16'h0000;
      ram[16'h003e] = 16'h0000;
      ram[16'h003f] = 16'h0000;
      ram[16'h0040] = 16'h0000;
      ram[16'h0041] = 16'h0000;
      ram[16'h0042] = 16'h0000;
      ram[16'h0043] = 16'h0000;
      ram[16'h0044] = 16'h0000;
      ram[16'h0045] = 16'h0000;
      ram[16'h0046] = 16'h0000;
      ram[16'h0047] = 16'h0000;
      ram[16'h0048] = 16'h0000;
      ram[16'h0049] = 16'h0000;
      ram[16'h004a] = 16'h0000;
      ram[16'h004b] = 16'h0000;
      ram[16'h004c] = 16'h0000;
      ram[16'h004d] = 16'h0000;
      ram[16'h004e] = 16'h0000;
      ram[16'h004f] = 16'h0000;
      ram[16'h0050] = 16'h0000;
      ram[16'h0051] = 16'h0000;
      ram[16'h0052] = 16'h0000;
      ram[16'h0053] = 16'h0000;
      ram[16'h0054] = 16'h0000;
      ram[16'h0055] = 16'h0000;
      ram[16'h0056] = 16'h0000;
      ram[16'h0057] = 16'h0000;
      ram[16'h0058] = 16'h0000;
      ram[16'h0059] = 16'h0000;
      ram[16'h005a] = 16'h0000;
      ram[16'h005b] = 16'h0000;
      ram[16'h005c] = 16'h0000;
      ram[16'h005d] = 16'h0000;
      ram[16'h005e] = 16'h0000;
      ram[16'h005f] = 16'h0000;
      ram[16'h0060] = 16'h0000;
      ram[16'h0061] = 16'h0000;
      ram[16'h0062] = 16'h0000;
      ram[16'h0063] = 16'h0000;
      ram[16'h0064] = 16'h0000;
      ram[16'h0065] = 16'h0000;
      ram[16'h0066] = 16'h0000;
      ram[16'h0067] = 16'h0000;
      ram[16'h0068] = 16'h0000;
      ram[16'h0069] = 16'h0000;
      ram[16'h006a] = 16'h0000;
      ram[16'h006b] = 16'h0000;
      ram[16'h006c] = 16'h0000;
      ram[16'h006d] = 16'h0000;
      ram[16'h006e] = 16'h0000;
      ram[16'h006f] = 16'h0000;
      ram[16'h0070] = 16'h0000;
      ram[16'h0071] = 16'h0000;
      ram[16'h0072] = 16'h0000;
      ram[16'h0073] = 16'h0000;
      ram[16'h0074] = 16'h0000;
      ram[16'h0075] = 16'h0000;
      ram[16'h0076] = 16'h0000;
      ram[16'h0077] = 16'h0000;
      ram[16'h0078] = 16'h0000;
      ram[16'h0079] = 16'h0000;
      ram[16'h007a] = 16'h0000;
      ram[16'h007b] = 16'h0000;
      ram[16'h007c] = 16'h0000;
      ram[16'h007d] = 16'h0000;
      ram[16'h007e] = 16'h0000;
      ram[16'h007f] = 16'h0000;
      ram[16'h0080] = 16'h0000;
      ram[16'h0081] = 16'h0000;
      ram[16'h0082] = 16'h0000;
      ram[16'h0083] = 16'h0000;
      ram[16'h0084] = 16'h0000;
      ram[16'h0085] = 16'h0000;
      ram[16'h0086] = 16'h0000;
      ram[16'h0087] = 16'h0000;
      ram[16'h0088] = 16'h0000;
      ram[16'h0089] = 16'h0000;
      ram[16'h008a] = 16'h0000;
      ram[16'h008b] = 16'h0000;
      ram[16'h008c] = 16'h0000;
      ram[16'h008d] = 16'h0000;
      ram[16'h008e] = 16'h0000;
      ram[16'h008f] = 16'h0000;
      ram[16'h0090] = 16'h0000;
      ram[16'h0091] = 16'h0000;
      ram[16'h0092] = 16'h0000;
      ram[16'h0093] = 16'h0000;
      ram[16'h0094] = 16'h0000;
      ram[16'h0095] = 16'h0000;
      ram[16'h0096] = 16'h0000;
      ram[16'h0097] = 16'h0000;
      ram[16'h0098] = 16'h0000;
      ram[16'h0099] = 16'h0000;
      ram[16'h009a] = 16'h0000;
      ram[16'h009b] = 16'h0000;
      ram[16'h009c] = 16'h0000;
      ram[16'h009d] = 16'h0000;
      ram[16'h009e] = 16'h0000;
      ram[16'h009f] = 16'h0000;
      ram[16'h00a0] = 16'h0000;
      ram[16'h00a1] = 16'h0000;
      ram[16'h00a2] = 16'h0000;
      ram[16'h00a3] = 16'h0000;
      ram[16'h00a4] = 16'h0000;
      ram[16'h00a5] = 16'h0000;
      ram[16'h00a6] = 16'h0000;
      ram[16'h00a7] = 16'h0000;
      ram[16'h00a8] = 16'h0000;
      ram[16'h00a9] = 16'h0000;
      ram[16'h00aa] = 16'h0000;
      ram[16'h00ab] = 16'h0000;
      ram[16'h00ac] = 16'h0000;
      ram[16'h00ad] = 16'h0000;
      ram[16'h00ae] = 16'h0000;
      ram[16'h00af] = 16'h0000;
      ram[16'h00b0] = 16'h0000;
      ram[16'h00b1] = 16'h0000;
      ram[16'h00b2] = 16'h0000;
      ram[16'h00b3] = 16'h0000;
      ram[16'h00b4] = 16'h0000;
      ram[16'h00b5] = 16'h0000;
      ram[16'h00b6] = 16'h0000;
      ram[16'h00b7] = 16'h0000;
      ram[16'h00b8] = 16'h0000;
      ram[16'h00b9] = 16'h0000;
      ram[16'h00ba] = 16'h0000;
      ram[16'h00bb] = 16'h0000;
      ram[16'h00bc] = 16'h0000;
      ram[16'h00bd] = 16'h0000;
      ram[16'h00be] = 16'h0000;
      ram[16'h00bf] = 16'h0000;
      ram[16'h00c0] = 16'h0000;
      ram[16'h00c1] = 16'h0000;
      ram[16'h00c2] = 16'h0000;
      ram[16'h00c3] = 16'h0000;
      ram[16'h00c4] = 16'h0000;
      ram[16'h00c5] = 16'h0000;
      ram[16'h00c6] = 16'h0000;
      ram[16'h00c7] = 16'h0000;
      ram[16'h00c8] = 16'h0000;
      ram[16'h00c9] = 16'h0000;
      ram[16'h00ca] = 16'h0000;
      ram[16'h00cb] = 16'h0000;
      ram[16'h00cc] = 16'h0000;
      ram[16'h00cd] = 16'h0000;
      ram[16'h00ce] = 16'h0000;
      ram[16'h00cf] = 16'h0000;
      ram[16'h00d0] = 16'h0000;
      ram[16'h00d1] = 16'h0000;
      ram[16'h00d2] = 16'h0000;
      ram[16'h00d3] = 16'h0000;
      ram[16'h00d4] = 16'h0000;
      ram[16'h00d5] = 16'h0000;
      ram[16'h00d6] = 16'h0000;
      ram[16'h00d7] = 16'h0000;
      ram[16'h00d8] = 16'h0000;
      ram[16'h00d9] = 16'h0000;
      ram[16'h00da] = 16'h0000;
      ram[16'h00db] = 16'h0000;
      ram[16'h00dc] = 16'h0000;
      ram[16'h00dd] = 16'h0000;
      ram[16'h00de] = 16'h0000;
      ram[16'h00df] = 16'h0000;
      ram[16'h00e0] = 16'h0000;
      ram[16'h00e1] = 16'h0000;
      ram[16'h00e2] = 16'h0000;
      ram[16'h00e3] = 16'h0000;
      ram[16'h00e4] = 16'h0000;
      ram[16'h00e5] = 16'h0000;
      ram[16'h00e6] = 16'h0000;
      ram[16'h00e7] = 16'h0000;
      ram[16'h00e8] = 16'h0000;
      ram[16'h00e9] = 16'h0000;
      ram[16'h00ea] = 16'h0000;
      ram[16'h00eb] = 16'h0000;
      ram[16'h00ec] = 16'h0000;
      ram[16'h00ed] = 16'h0000;
      ram[16'h00ee] = 16'h0000;
      ram[16'h00ef] = 16'h0000;
      ram[16'h00f0] = 16'h0000;
      ram[16'h00f1] = 16'h0000;
      ram[16'h00f2] = 16'h0000;
      ram[16'h00f3] = 16'h0000;
      ram[16'h00f4] = 16'h0000;
      ram[16'h00f5] = 16'h0000;
      ram[16'h00f6] = 16'h0000;
      ram[16'h00f7] = 16'h0000;
      ram[16'h00f8] = 16'h0000;
      ram[16'h00f9] = 16'h0000;
      ram[16'h00fa] = 16'h0000;
      ram[16'h00fb] = 16'h0000;
      ram[16'h00fc] = 16'h0000;
      ram[16'h00fd] = 16'h0000;
      ram[16'h00fe] = 16'h0000;
      ram[16'h00ff] = 16'h0000;
    end

endmodule
